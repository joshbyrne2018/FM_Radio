library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


package CoArray_pkg is

     type CoArray is array (integer range <>) of integer;

end package CoArray_pkg;